VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RF
  CLASS BLOCK ;
  FOREIGN RF ;
  ORIGIN 0.000 0.000 ;
  SIZE 590.000 BY 820.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.720 4.000 800.320 ;
    END
  END clk
  PIN raddr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 10.240 590.000 10.840 ;
    END
  END raddr0[0]
  PIN raddr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 146.240 590.000 146.840 ;
    END
  END raddr0[1]
  PIN raddr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 282.240 590.000 282.840 ;
    END
  END raddr0[2]
  PIN raddr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 418.240 590.000 418.840 ;
    END
  END raddr0[3]
  PIN raddr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 554.240 590.000 554.840 ;
    END
  END raddr0[4]
  PIN raddr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 690.240 590.000 690.840 ;
    END
  END raddr0[5]
  PIN raddr1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 27.240 590.000 27.840 ;
    END
  END raddr1[0]
  PIN raddr1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 163.240 590.000 163.840 ;
    END
  END raddr1[1]
  PIN raddr1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 299.240 590.000 299.840 ;
    END
  END raddr1[2]
  PIN raddr1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 435.240 590.000 435.840 ;
    END
  END raddr1[3]
  PIN raddr1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 571.240 590.000 571.840 ;
    END
  END raddr1[4]
  PIN raddr1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 707.240 590.000 707.840 ;
    END
  END raddr1[5]
  PIN raddr2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 44.240 590.000 44.840 ;
    END
  END raddr2[0]
  PIN raddr2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 180.240 590.000 180.840 ;
    END
  END raddr2[1]
  PIN raddr2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 316.240 590.000 316.840 ;
    END
  END raddr2[2]
  PIN raddr2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 452.240 590.000 452.840 ;
    END
  END raddr2[3]
  PIN raddr2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 588.240 590.000 588.840 ;
    END
  END raddr2[4]
  PIN raddr2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 724.240 590.000 724.840 ;
    END
  END raddr2[5]
  PIN raddr3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 61.240 590.000 61.840 ;
    END
  END raddr3[0]
  PIN raddr3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 197.240 590.000 197.840 ;
    END
  END raddr3[1]
  PIN raddr3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 333.240 590.000 333.840 ;
    END
  END raddr3[2]
  PIN raddr3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 469.240 590.000 469.840 ;
    END
  END raddr3[3]
  PIN raddr3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 605.240 590.000 605.840 ;
    END
  END raddr3[4]
  PIN raddr3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 741.240 590.000 741.840 ;
    END
  END raddr3[5]
  PIN raddr4[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 78.240 590.000 78.840 ;
    END
  END raddr4[0]
  PIN raddr4[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 214.240 590.000 214.840 ;
    END
  END raddr4[1]
  PIN raddr4[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 350.240 590.000 350.840 ;
    END
  END raddr4[2]
  PIN raddr4[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 486.240 590.000 486.840 ;
    END
  END raddr4[3]
  PIN raddr4[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 622.240 590.000 622.840 ;
    END
  END raddr4[4]
  PIN raddr4[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 758.240 590.000 758.840 ;
    END
  END raddr4[5]
  PIN raddr5[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 95.240 590.000 95.840 ;
    END
  END raddr5[0]
  PIN raddr5[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 231.240 590.000 231.840 ;
    END
  END raddr5[1]
  PIN raddr5[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 367.240 590.000 367.840 ;
    END
  END raddr5[2]
  PIN raddr5[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 503.240 590.000 503.840 ;
    END
  END raddr5[3]
  PIN raddr5[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 639.240 590.000 639.840 ;
    END
  END raddr5[4]
  PIN raddr5[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 775.240 590.000 775.840 ;
    END
  END raddr5[5]
  PIN raddr6[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 112.240 590.000 112.840 ;
    END
  END raddr6[0]
  PIN raddr6[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 248.240 590.000 248.840 ;
    END
  END raddr6[1]
  PIN raddr6[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 384.240 590.000 384.840 ;
    END
  END raddr6[2]
  PIN raddr6[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 520.240 590.000 520.840 ;
    END
  END raddr6[3]
  PIN raddr6[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 656.240 590.000 656.840 ;
    END
  END raddr6[4]
  PIN raddr6[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 792.240 590.000 792.840 ;
    END
  END raddr6[5]
  PIN raddr7[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 129.240 590.000 129.840 ;
    END
  END raddr7[0]
  PIN raddr7[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 265.240 590.000 265.840 ;
    END
  END raddr7[1]
  PIN raddr7[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 401.240 590.000 401.840 ;
    END
  END raddr7[2]
  PIN raddr7[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 537.240 590.000 537.840 ;
    END
  END raddr7[3]
  PIN raddr7[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 673.240 590.000 673.840 ;
    END
  END raddr7[4]
  PIN raddr7[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.000 809.240 590.000 809.840 ;
    END
  END raddr7[5]
  PIN rdata0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END rdata0[0]
  PIN rdata0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END rdata0[10]
  PIN rdata0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END rdata0[11]
  PIN rdata0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END rdata0[12]
  PIN rdata0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END rdata0[13]
  PIN rdata0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END rdata0[14]
  PIN rdata0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 4.000 ;
    END
  END rdata0[15]
  PIN rdata0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END rdata0[16]
  PIN rdata0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END rdata0[17]
  PIN rdata0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END rdata0[18]
  PIN rdata0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END rdata0[19]
  PIN rdata0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END rdata0[1]
  PIN rdata0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END rdata0[20]
  PIN rdata0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END rdata0[21]
  PIN rdata0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END rdata0[22]
  PIN rdata0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END rdata0[23]
  PIN rdata0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END rdata0[24]
  PIN rdata0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END rdata0[25]
  PIN rdata0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END rdata0[26]
  PIN rdata0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 0.000 498.550 4.000 ;
    END
  END rdata0[27]
  PIN rdata0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 0.000 516.950 4.000 ;
    END
  END rdata0[28]
  PIN rdata0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 0.000 535.350 4.000 ;
    END
  END rdata0[29]
  PIN rdata0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END rdata0[2]
  PIN rdata0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END rdata0[30]
  PIN rdata0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 0.000 572.150 4.000 ;
    END
  END rdata0[31]
  PIN rdata0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END rdata0[3]
  PIN rdata0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END rdata0[4]
  PIN rdata0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END rdata0[5]
  PIN rdata0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END rdata0[6]
  PIN rdata0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END rdata0[7]
  PIN rdata0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END rdata0[8]
  PIN rdata0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END rdata0[9]
  PIN rdata1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END rdata1[0]
  PIN rdata1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END rdata1[10]
  PIN rdata1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END rdata1[11]
  PIN rdata1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END rdata1[12]
  PIN rdata1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END rdata1[13]
  PIN rdata1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END rdata1[14]
  PIN rdata1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END rdata1[15]
  PIN rdata1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END rdata1[16]
  PIN rdata1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END rdata1[17]
  PIN rdata1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END rdata1[18]
  PIN rdata1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END rdata1[19]
  PIN rdata1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END rdata1[1]
  PIN rdata1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END rdata1[20]
  PIN rdata1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END rdata1[21]
  PIN rdata1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END rdata1[22]
  PIN rdata1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 4.000 ;
    END
  END rdata1[23]
  PIN rdata1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 0.000 445.650 4.000 ;
    END
  END rdata1[24]
  PIN rdata1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END rdata1[25]
  PIN rdata1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END rdata1[26]
  PIN rdata1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END rdata1[27]
  PIN rdata1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 0.000 519.250 4.000 ;
    END
  END rdata1[28]
  PIN rdata1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END rdata1[29]
  PIN rdata1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END rdata1[2]
  PIN rdata1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 0.000 556.050 4.000 ;
    END
  END rdata1[30]
  PIN rdata1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END rdata1[31]
  PIN rdata1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END rdata1[3]
  PIN rdata1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END rdata1[4]
  PIN rdata1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END rdata1[5]
  PIN rdata1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END rdata1[6]
  PIN rdata1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END rdata1[7]
  PIN rdata1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END rdata1[8]
  PIN rdata1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END rdata1[9]
  PIN rdata2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END rdata2[0]
  PIN rdata2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END rdata2[10]
  PIN rdata2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END rdata2[11]
  PIN rdata2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 0.000 227.150 4.000 ;
    END
  END rdata2[12]
  PIN rdata2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END rdata2[13]
  PIN rdata2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END rdata2[14]
  PIN rdata2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END rdata2[15]
  PIN rdata2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END rdata2[16]
  PIN rdata2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END rdata2[17]
  PIN rdata2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END rdata2[18]
  PIN rdata2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 4.000 ;
    END
  END rdata2[19]
  PIN rdata2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END rdata2[1]
  PIN rdata2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END rdata2[20]
  PIN rdata2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END rdata2[21]
  PIN rdata2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 4.000 ;
    END
  END rdata2[22]
  PIN rdata2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END rdata2[23]
  PIN rdata2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END rdata2[24]
  PIN rdata2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 0.000 466.350 4.000 ;
    END
  END rdata2[25]
  PIN rdata2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 0.000 484.750 4.000 ;
    END
  END rdata2[26]
  PIN rdata2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 0.000 503.150 4.000 ;
    END
  END rdata2[27]
  PIN rdata2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END rdata2[28]
  PIN rdata2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END rdata2[29]
  PIN rdata2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END rdata2[2]
  PIN rdata2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 0.000 558.350 4.000 ;
    END
  END rdata2[30]
  PIN rdata2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END rdata2[31]
  PIN rdata2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END rdata2[3]
  PIN rdata2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END rdata2[4]
  PIN rdata2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END rdata2[5]
  PIN rdata2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END rdata2[6]
  PIN rdata2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END rdata2[7]
  PIN rdata2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END rdata2[8]
  PIN rdata2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END rdata2[9]
  PIN rdata3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END rdata3[0]
  PIN rdata3[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END rdata3[10]
  PIN rdata3[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END rdata3[11]
  PIN rdata3[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END rdata3[12]
  PIN rdata3[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END rdata3[13]
  PIN rdata3[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END rdata3[14]
  PIN rdata3[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END rdata3[15]
  PIN rdata3[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END rdata3[16]
  PIN rdata3[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END rdata3[17]
  PIN rdata3[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END rdata3[18]
  PIN rdata3[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END rdata3[19]
  PIN rdata3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END rdata3[1]
  PIN rdata3[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END rdata3[20]
  PIN rdata3[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END rdata3[21]
  PIN rdata3[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END rdata3[22]
  PIN rdata3[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END rdata3[23]
  PIN rdata3[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END rdata3[24]
  PIN rdata3[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END rdata3[25]
  PIN rdata3[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 4.000 ;
    END
  END rdata3[26]
  PIN rdata3[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END rdata3[27]
  PIN rdata3[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 0.000 523.850 4.000 ;
    END
  END rdata3[28]
  PIN rdata3[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.970 0.000 542.250 4.000 ;
    END
  END rdata3[29]
  PIN rdata3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END rdata3[2]
  PIN rdata3[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END rdata3[30]
  PIN rdata3[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.770 0.000 579.050 4.000 ;
    END
  END rdata3[31]
  PIN rdata3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END rdata3[3]
  PIN rdata3[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END rdata3[4]
  PIN rdata3[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END rdata3[5]
  PIN rdata3[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END rdata3[6]
  PIN rdata3[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END rdata3[7]
  PIN rdata3[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END rdata3[8]
  PIN rdata3[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END rdata3[9]
  PIN rdata4[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END rdata4[0]
  PIN rdata4[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END rdata4[10]
  PIN rdata4[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END rdata4[11]
  PIN rdata4[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END rdata4[12]
  PIN rdata4[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END rdata4[13]
  PIN rdata4[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END rdata4[14]
  PIN rdata4[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END rdata4[15]
  PIN rdata4[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END rdata4[16]
  PIN rdata4[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END rdata4[17]
  PIN rdata4[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END rdata4[18]
  PIN rdata4[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END rdata4[19]
  PIN rdata4[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END rdata4[1]
  PIN rdata4[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END rdata4[20]
  PIN rdata4[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END rdata4[21]
  PIN rdata4[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END rdata4[22]
  PIN rdata4[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 0.000 434.150 4.000 ;
    END
  END rdata4[23]
  PIN rdata4[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END rdata4[24]
  PIN rdata4[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 4.000 ;
    END
  END rdata4[25]
  PIN rdata4[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END rdata4[26]
  PIN rdata4[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END rdata4[27]
  PIN rdata4[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 0.000 526.150 4.000 ;
    END
  END rdata4[28]
  PIN rdata4[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END rdata4[29]
  PIN rdata4[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END rdata4[2]
  PIN rdata4[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END rdata4[30]
  PIN rdata4[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END rdata4[31]
  PIN rdata4[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END rdata4[3]
  PIN rdata4[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END rdata4[4]
  PIN rdata4[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END rdata4[5]
  PIN rdata4[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END rdata4[6]
  PIN rdata4[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END rdata4[7]
  PIN rdata4[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END rdata4[8]
  PIN rdata4[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END rdata4[9]
  PIN rdata5[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END rdata5[0]
  PIN rdata5[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END rdata5[10]
  PIN rdata5[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END rdata5[11]
  PIN rdata5[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END rdata5[12]
  PIN rdata5[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END rdata5[13]
  PIN rdata5[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END rdata5[14]
  PIN rdata5[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END rdata5[15]
  PIN rdata5[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END rdata5[16]
  PIN rdata5[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END rdata5[17]
  PIN rdata5[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END rdata5[18]
  PIN rdata5[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END rdata5[19]
  PIN rdata5[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END rdata5[1]
  PIN rdata5[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END rdata5[20]
  PIN rdata5[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END rdata5[21]
  PIN rdata5[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END rdata5[22]
  PIN rdata5[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END rdata5[23]
  PIN rdata5[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 0.000 454.850 4.000 ;
    END
  END rdata5[24]
  PIN rdata5[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 0.000 473.250 4.000 ;
    END
  END rdata5[25]
  PIN rdata5[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END rdata5[26]
  PIN rdata5[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 0.000 510.050 4.000 ;
    END
  END rdata5[27]
  PIN rdata5[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END rdata5[28]
  PIN rdata5[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 4.000 ;
    END
  END rdata5[29]
  PIN rdata5[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END rdata5[2]
  PIN rdata5[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END rdata5[30]
  PIN rdata5[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 0.000 583.650 4.000 ;
    END
  END rdata5[31]
  PIN rdata5[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END rdata5[3]
  PIN rdata5[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END rdata5[4]
  PIN rdata5[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END rdata5[5]
  PIN rdata5[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END rdata5[6]
  PIN rdata5[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END rdata5[7]
  PIN rdata5[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END rdata5[8]
  PIN rdata5[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END rdata5[9]
  PIN rdata6[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END rdata6[0]
  PIN rdata6[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END rdata6[10]
  PIN rdata6[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END rdata6[11]
  PIN rdata6[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END rdata6[12]
  PIN rdata6[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END rdata6[13]
  PIN rdata6[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END rdata6[14]
  PIN rdata6[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END rdata6[15]
  PIN rdata6[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END rdata6[16]
  PIN rdata6[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END rdata6[17]
  PIN rdata6[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END rdata6[18]
  PIN rdata6[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 0.000 365.150 4.000 ;
    END
  END rdata6[19]
  PIN rdata6[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END rdata6[1]
  PIN rdata6[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END rdata6[20]
  PIN rdata6[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 0.000 401.950 4.000 ;
    END
  END rdata6[21]
  PIN rdata6[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 0.000 420.350 4.000 ;
    END
  END rdata6[22]
  PIN rdata6[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END rdata6[23]
  PIN rdata6[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 0.000 457.150 4.000 ;
    END
  END rdata6[24]
  PIN rdata6[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END rdata6[25]
  PIN rdata6[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 0.000 493.950 4.000 ;
    END
  END rdata6[26]
  PIN rdata6[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END rdata6[27]
  PIN rdata6[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 0.000 530.750 4.000 ;
    END
  END rdata6[28]
  PIN rdata6[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 0.000 549.150 4.000 ;
    END
  END rdata6[29]
  PIN rdata6[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END rdata6[2]
  PIN rdata6[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 0.000 567.550 4.000 ;
    END
  END rdata6[30]
  PIN rdata6[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 4.000 ;
    END
  END rdata6[31]
  PIN rdata6[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END rdata6[3]
  PIN rdata6[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END rdata6[4]
  PIN rdata6[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END rdata6[5]
  PIN rdata6[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END rdata6[6]
  PIN rdata6[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END rdata6[7]
  PIN rdata6[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END rdata6[8]
  PIN rdata6[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END rdata6[9]
  PIN rdata7[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END rdata7[0]
  PIN rdata7[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END rdata7[10]
  PIN rdata7[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END rdata7[11]
  PIN rdata7[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END rdata7[12]
  PIN rdata7[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END rdata7[13]
  PIN rdata7[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END rdata7[14]
  PIN rdata7[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END rdata7[15]
  PIN rdata7[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END rdata7[16]
  PIN rdata7[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END rdata7[17]
  PIN rdata7[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END rdata7[18]
  PIN rdata7[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END rdata7[19]
  PIN rdata7[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END rdata7[1]
  PIN rdata7[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END rdata7[20]
  PIN rdata7[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 0.000 404.250 4.000 ;
    END
  END rdata7[21]
  PIN rdata7[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END rdata7[22]
  PIN rdata7[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END rdata7[23]
  PIN rdata7[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END rdata7[24]
  PIN rdata7[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 0.000 477.850 4.000 ;
    END
  END rdata7[25]
  PIN rdata7[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END rdata7[26]
  PIN rdata7[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 0.000 514.650 4.000 ;
    END
  END rdata7[27]
  PIN rdata7[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 0.000 533.050 4.000 ;
    END
  END rdata7[28]
  PIN rdata7[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END rdata7[29]
  PIN rdata7[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END rdata7[2]
  PIN rdata7[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 0.000 569.850 4.000 ;
    END
  END rdata7[30]
  PIN rdata7[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 4.000 ;
    END
  END rdata7[31]
  PIN rdata7[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END rdata7[3]
  PIN rdata7[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END rdata7[4]
  PIN rdata7[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END rdata7[5]
  PIN rdata7[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END rdata7[6]
  PIN rdata7[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END rdata7[7]
  PIN rdata7[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END rdata7[8]
  PIN rdata7[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END rdata7[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 808.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 808.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 808.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 808.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 808.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 808.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 808.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 808.080 ;
    END
  END vssd1
  PIN waddr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END waddr0[0]
  PIN waddr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END waddr0[1]
  PIN waddr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END waddr0[2]
  PIN waddr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END waddr0[3]
  PIN waddr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END waddr0[4]
  PIN waddr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.680 4.000 577.280 ;
    END
  END waddr0[5]
  PIN waddr1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END waddr1[0]
  PIN waddr1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END waddr1[1]
  PIN waddr1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END waddr1[2]
  PIN waddr1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END waddr1[3]
  PIN waddr1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END waddr1[4]
  PIN waddr1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 604.560 4.000 605.160 ;
    END
  END waddr1[5]
  PIN waddr2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END waddr2[0]
  PIN waddr2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END waddr2[1]
  PIN waddr2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END waddr2[2]
  PIN waddr2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END waddr2[3]
  PIN waddr2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END waddr2[4]
  PIN waddr2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END waddr2[5]
  PIN waddr3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END waddr3[0]
  PIN waddr3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END waddr3[1]
  PIN waddr3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END waddr3[2]
  PIN waddr3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.280 4.000 437.880 ;
    END
  END waddr3[3]
  PIN waddr3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.800 4.000 549.400 ;
    END
  END waddr3[4]
  PIN waddr3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END waddr3[5]
  PIN wdata0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 816.000 2.670 820.000 ;
    END
  END wdata0[0]
  PIN wdata0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 816.000 186.670 820.000 ;
    END
  END wdata0[10]
  PIN wdata0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 816.000 205.070 820.000 ;
    END
  END wdata0[11]
  PIN wdata0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 816.000 223.470 820.000 ;
    END
  END wdata0[12]
  PIN wdata0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 816.000 241.870 820.000 ;
    END
  END wdata0[13]
  PIN wdata0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 816.000 260.270 820.000 ;
    END
  END wdata0[14]
  PIN wdata0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 816.000 278.670 820.000 ;
    END
  END wdata0[15]
  PIN wdata0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 816.000 297.070 820.000 ;
    END
  END wdata0[16]
  PIN wdata0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 816.000 315.470 820.000 ;
    END
  END wdata0[17]
  PIN wdata0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 816.000 333.870 820.000 ;
    END
  END wdata0[18]
  PIN wdata0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 816.000 352.270 820.000 ;
    END
  END wdata0[19]
  PIN wdata0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 816.000 21.070 820.000 ;
    END
  END wdata0[1]
  PIN wdata0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 816.000 370.670 820.000 ;
    END
  END wdata0[20]
  PIN wdata0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 816.000 389.070 820.000 ;
    END
  END wdata0[21]
  PIN wdata0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 816.000 407.470 820.000 ;
    END
  END wdata0[22]
  PIN wdata0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 816.000 425.870 820.000 ;
    END
  END wdata0[23]
  PIN wdata0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 816.000 444.270 820.000 ;
    END
  END wdata0[24]
  PIN wdata0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 816.000 462.670 820.000 ;
    END
  END wdata0[25]
  PIN wdata0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 816.000 481.070 820.000 ;
    END
  END wdata0[26]
  PIN wdata0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 816.000 499.470 820.000 ;
    END
  END wdata0[27]
  PIN wdata0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 816.000 517.870 820.000 ;
    END
  END wdata0[28]
  PIN wdata0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 816.000 536.270 820.000 ;
    END
  END wdata0[29]
  PIN wdata0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 816.000 39.470 820.000 ;
    END
  END wdata0[2]
  PIN wdata0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 816.000 554.670 820.000 ;
    END
  END wdata0[30]
  PIN wdata0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 816.000 573.070 820.000 ;
    END
  END wdata0[31]
  PIN wdata0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 816.000 57.870 820.000 ;
    END
  END wdata0[3]
  PIN wdata0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 816.000 76.270 820.000 ;
    END
  END wdata0[4]
  PIN wdata0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 816.000 94.670 820.000 ;
    END
  END wdata0[5]
  PIN wdata0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 816.000 113.070 820.000 ;
    END
  END wdata0[6]
  PIN wdata0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 816.000 131.470 820.000 ;
    END
  END wdata0[7]
  PIN wdata0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 816.000 149.870 820.000 ;
    END
  END wdata0[8]
  PIN wdata0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 816.000 168.270 820.000 ;
    END
  END wdata0[9]
  PIN wdata1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 816.000 7.270 820.000 ;
    END
  END wdata1[0]
  PIN wdata1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 816.000 191.270 820.000 ;
    END
  END wdata1[10]
  PIN wdata1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 816.000 209.670 820.000 ;
    END
  END wdata1[11]
  PIN wdata1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 816.000 228.070 820.000 ;
    END
  END wdata1[12]
  PIN wdata1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 816.000 246.470 820.000 ;
    END
  END wdata1[13]
  PIN wdata1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 816.000 264.870 820.000 ;
    END
  END wdata1[14]
  PIN wdata1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 816.000 283.270 820.000 ;
    END
  END wdata1[15]
  PIN wdata1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 816.000 301.670 820.000 ;
    END
  END wdata1[16]
  PIN wdata1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 816.000 320.070 820.000 ;
    END
  END wdata1[17]
  PIN wdata1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 816.000 338.470 820.000 ;
    END
  END wdata1[18]
  PIN wdata1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 816.000 356.870 820.000 ;
    END
  END wdata1[19]
  PIN wdata1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 816.000 25.670 820.000 ;
    END
  END wdata1[1]
  PIN wdata1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 816.000 375.270 820.000 ;
    END
  END wdata1[20]
  PIN wdata1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 816.000 393.670 820.000 ;
    END
  END wdata1[21]
  PIN wdata1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 816.000 412.070 820.000 ;
    END
  END wdata1[22]
  PIN wdata1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 816.000 430.470 820.000 ;
    END
  END wdata1[23]
  PIN wdata1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 816.000 448.870 820.000 ;
    END
  END wdata1[24]
  PIN wdata1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 816.000 467.270 820.000 ;
    END
  END wdata1[25]
  PIN wdata1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 816.000 485.670 820.000 ;
    END
  END wdata1[26]
  PIN wdata1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 816.000 504.070 820.000 ;
    END
  END wdata1[27]
  PIN wdata1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 816.000 522.470 820.000 ;
    END
  END wdata1[28]
  PIN wdata1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 816.000 540.870 820.000 ;
    END
  END wdata1[29]
  PIN wdata1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 816.000 44.070 820.000 ;
    END
  END wdata1[2]
  PIN wdata1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 816.000 559.270 820.000 ;
    END
  END wdata1[30]
  PIN wdata1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 816.000 577.670 820.000 ;
    END
  END wdata1[31]
  PIN wdata1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 816.000 62.470 820.000 ;
    END
  END wdata1[3]
  PIN wdata1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 816.000 80.870 820.000 ;
    END
  END wdata1[4]
  PIN wdata1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 816.000 99.270 820.000 ;
    END
  END wdata1[5]
  PIN wdata1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 816.000 117.670 820.000 ;
    END
  END wdata1[6]
  PIN wdata1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 816.000 136.070 820.000 ;
    END
  END wdata1[7]
  PIN wdata1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 816.000 154.470 820.000 ;
    END
  END wdata1[8]
  PIN wdata1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 816.000 172.870 820.000 ;
    END
  END wdata1[9]
  PIN wdata2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 816.000 11.870 820.000 ;
    END
  END wdata2[0]
  PIN wdata2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 816.000 195.870 820.000 ;
    END
  END wdata2[10]
  PIN wdata2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 816.000 214.270 820.000 ;
    END
  END wdata2[11]
  PIN wdata2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 816.000 232.670 820.000 ;
    END
  END wdata2[12]
  PIN wdata2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 816.000 251.070 820.000 ;
    END
  END wdata2[13]
  PIN wdata2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 816.000 269.470 820.000 ;
    END
  END wdata2[14]
  PIN wdata2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 816.000 287.870 820.000 ;
    END
  END wdata2[15]
  PIN wdata2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 816.000 306.270 820.000 ;
    END
  END wdata2[16]
  PIN wdata2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 816.000 324.670 820.000 ;
    END
  END wdata2[17]
  PIN wdata2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 816.000 343.070 820.000 ;
    END
  END wdata2[18]
  PIN wdata2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 816.000 361.470 820.000 ;
    END
  END wdata2[19]
  PIN wdata2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 816.000 30.270 820.000 ;
    END
  END wdata2[1]
  PIN wdata2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 816.000 379.870 820.000 ;
    END
  END wdata2[20]
  PIN wdata2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 816.000 398.270 820.000 ;
    END
  END wdata2[21]
  PIN wdata2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 816.000 416.670 820.000 ;
    END
  END wdata2[22]
  PIN wdata2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 816.000 435.070 820.000 ;
    END
  END wdata2[23]
  PIN wdata2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 816.000 453.470 820.000 ;
    END
  END wdata2[24]
  PIN wdata2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 816.000 471.870 820.000 ;
    END
  END wdata2[25]
  PIN wdata2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 816.000 490.270 820.000 ;
    END
  END wdata2[26]
  PIN wdata2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 816.000 508.670 820.000 ;
    END
  END wdata2[27]
  PIN wdata2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 816.000 527.070 820.000 ;
    END
  END wdata2[28]
  PIN wdata2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 816.000 545.470 820.000 ;
    END
  END wdata2[29]
  PIN wdata2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 816.000 48.670 820.000 ;
    END
  END wdata2[2]
  PIN wdata2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 816.000 563.870 820.000 ;
    END
  END wdata2[30]
  PIN wdata2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 816.000 582.270 820.000 ;
    END
  END wdata2[31]
  PIN wdata2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 816.000 67.070 820.000 ;
    END
  END wdata2[3]
  PIN wdata2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 816.000 85.470 820.000 ;
    END
  END wdata2[4]
  PIN wdata2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 816.000 103.870 820.000 ;
    END
  END wdata2[5]
  PIN wdata2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 816.000 122.270 820.000 ;
    END
  END wdata2[6]
  PIN wdata2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 816.000 140.670 820.000 ;
    END
  END wdata2[7]
  PIN wdata2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 816.000 159.070 820.000 ;
    END
  END wdata2[8]
  PIN wdata2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 816.000 177.470 820.000 ;
    END
  END wdata2[9]
  PIN wdata3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 816.000 16.470 820.000 ;
    END
  END wdata3[0]
  PIN wdata3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 816.000 200.470 820.000 ;
    END
  END wdata3[10]
  PIN wdata3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 816.000 218.870 820.000 ;
    END
  END wdata3[11]
  PIN wdata3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 816.000 237.270 820.000 ;
    END
  END wdata3[12]
  PIN wdata3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 816.000 255.670 820.000 ;
    END
  END wdata3[13]
  PIN wdata3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 816.000 274.070 820.000 ;
    END
  END wdata3[14]
  PIN wdata3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 816.000 292.470 820.000 ;
    END
  END wdata3[15]
  PIN wdata3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 816.000 310.870 820.000 ;
    END
  END wdata3[16]
  PIN wdata3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 816.000 329.270 820.000 ;
    END
  END wdata3[17]
  PIN wdata3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 816.000 347.670 820.000 ;
    END
  END wdata3[18]
  PIN wdata3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 816.000 366.070 820.000 ;
    END
  END wdata3[19]
  PIN wdata3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 816.000 34.870 820.000 ;
    END
  END wdata3[1]
  PIN wdata3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 816.000 384.470 820.000 ;
    END
  END wdata3[20]
  PIN wdata3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 816.000 402.870 820.000 ;
    END
  END wdata3[21]
  PIN wdata3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 816.000 421.270 820.000 ;
    END
  END wdata3[22]
  PIN wdata3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 816.000 439.670 820.000 ;
    END
  END wdata3[23]
  PIN wdata3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 816.000 458.070 820.000 ;
    END
  END wdata3[24]
  PIN wdata3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 816.000 476.470 820.000 ;
    END
  END wdata3[25]
  PIN wdata3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 816.000 494.870 820.000 ;
    END
  END wdata3[26]
  PIN wdata3[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 816.000 513.270 820.000 ;
    END
  END wdata3[27]
  PIN wdata3[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 816.000 531.670 820.000 ;
    END
  END wdata3[28]
  PIN wdata3[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 816.000 550.070 820.000 ;
    END
  END wdata3[29]
  PIN wdata3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 816.000 53.270 820.000 ;
    END
  END wdata3[2]
  PIN wdata3[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 816.000 568.470 820.000 ;
    END
  END wdata3[30]
  PIN wdata3[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 816.000 586.870 820.000 ;
    END
  END wdata3[31]
  PIN wdata3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 816.000 71.670 820.000 ;
    END
  END wdata3[3]
  PIN wdata3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 816.000 90.070 820.000 ;
    END
  END wdata3[4]
  PIN wdata3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 816.000 108.470 820.000 ;
    END
  END wdata3[5]
  PIN wdata3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 816.000 126.870 820.000 ;
    END
  END wdata3[6]
  PIN wdata3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 816.000 145.270 820.000 ;
    END
  END wdata3[7]
  PIN wdata3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 816.000 163.670 820.000 ;
    END
  END wdata3[8]
  PIN wdata3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 816.000 182.070 820.000 ;
    END
  END wdata3[9]
  PIN wen0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END wen0
  PIN wen1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.080 4.000 716.680 ;
    END
  END wen1
  PIN wen2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END wen2
  PIN wen3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END wen3
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 584.200 807.925 ;
      LAYER met1 ;
        RECT 1.450 4.460 589.650 808.080 ;
      LAYER met2 ;
        RECT 1.480 815.720 2.110 816.410 ;
        RECT 2.950 815.720 6.710 816.410 ;
        RECT 7.550 815.720 11.310 816.410 ;
        RECT 12.150 815.720 15.910 816.410 ;
        RECT 16.750 815.720 20.510 816.410 ;
        RECT 21.350 815.720 25.110 816.410 ;
        RECT 25.950 815.720 29.710 816.410 ;
        RECT 30.550 815.720 34.310 816.410 ;
        RECT 35.150 815.720 38.910 816.410 ;
        RECT 39.750 815.720 43.510 816.410 ;
        RECT 44.350 815.720 48.110 816.410 ;
        RECT 48.950 815.720 52.710 816.410 ;
        RECT 53.550 815.720 57.310 816.410 ;
        RECT 58.150 815.720 61.910 816.410 ;
        RECT 62.750 815.720 66.510 816.410 ;
        RECT 67.350 815.720 71.110 816.410 ;
        RECT 71.950 815.720 75.710 816.410 ;
        RECT 76.550 815.720 80.310 816.410 ;
        RECT 81.150 815.720 84.910 816.410 ;
        RECT 85.750 815.720 89.510 816.410 ;
        RECT 90.350 815.720 94.110 816.410 ;
        RECT 94.950 815.720 98.710 816.410 ;
        RECT 99.550 815.720 103.310 816.410 ;
        RECT 104.150 815.720 107.910 816.410 ;
        RECT 108.750 815.720 112.510 816.410 ;
        RECT 113.350 815.720 117.110 816.410 ;
        RECT 117.950 815.720 121.710 816.410 ;
        RECT 122.550 815.720 126.310 816.410 ;
        RECT 127.150 815.720 130.910 816.410 ;
        RECT 131.750 815.720 135.510 816.410 ;
        RECT 136.350 815.720 140.110 816.410 ;
        RECT 140.950 815.720 144.710 816.410 ;
        RECT 145.550 815.720 149.310 816.410 ;
        RECT 150.150 815.720 153.910 816.410 ;
        RECT 154.750 815.720 158.510 816.410 ;
        RECT 159.350 815.720 163.110 816.410 ;
        RECT 163.950 815.720 167.710 816.410 ;
        RECT 168.550 815.720 172.310 816.410 ;
        RECT 173.150 815.720 176.910 816.410 ;
        RECT 177.750 815.720 181.510 816.410 ;
        RECT 182.350 815.720 186.110 816.410 ;
        RECT 186.950 815.720 190.710 816.410 ;
        RECT 191.550 815.720 195.310 816.410 ;
        RECT 196.150 815.720 199.910 816.410 ;
        RECT 200.750 815.720 204.510 816.410 ;
        RECT 205.350 815.720 209.110 816.410 ;
        RECT 209.950 815.720 213.710 816.410 ;
        RECT 214.550 815.720 218.310 816.410 ;
        RECT 219.150 815.720 222.910 816.410 ;
        RECT 223.750 815.720 227.510 816.410 ;
        RECT 228.350 815.720 232.110 816.410 ;
        RECT 232.950 815.720 236.710 816.410 ;
        RECT 237.550 815.720 241.310 816.410 ;
        RECT 242.150 815.720 245.910 816.410 ;
        RECT 246.750 815.720 250.510 816.410 ;
        RECT 251.350 815.720 255.110 816.410 ;
        RECT 255.950 815.720 259.710 816.410 ;
        RECT 260.550 815.720 264.310 816.410 ;
        RECT 265.150 815.720 268.910 816.410 ;
        RECT 269.750 815.720 273.510 816.410 ;
        RECT 274.350 815.720 278.110 816.410 ;
        RECT 278.950 815.720 282.710 816.410 ;
        RECT 283.550 815.720 287.310 816.410 ;
        RECT 288.150 815.720 291.910 816.410 ;
        RECT 292.750 815.720 296.510 816.410 ;
        RECT 297.350 815.720 301.110 816.410 ;
        RECT 301.950 815.720 305.710 816.410 ;
        RECT 306.550 815.720 310.310 816.410 ;
        RECT 311.150 815.720 314.910 816.410 ;
        RECT 315.750 815.720 319.510 816.410 ;
        RECT 320.350 815.720 324.110 816.410 ;
        RECT 324.950 815.720 328.710 816.410 ;
        RECT 329.550 815.720 333.310 816.410 ;
        RECT 334.150 815.720 337.910 816.410 ;
        RECT 338.750 815.720 342.510 816.410 ;
        RECT 343.350 815.720 347.110 816.410 ;
        RECT 347.950 815.720 351.710 816.410 ;
        RECT 352.550 815.720 356.310 816.410 ;
        RECT 357.150 815.720 360.910 816.410 ;
        RECT 361.750 815.720 365.510 816.410 ;
        RECT 366.350 815.720 370.110 816.410 ;
        RECT 370.950 815.720 374.710 816.410 ;
        RECT 375.550 815.720 379.310 816.410 ;
        RECT 380.150 815.720 383.910 816.410 ;
        RECT 384.750 815.720 388.510 816.410 ;
        RECT 389.350 815.720 393.110 816.410 ;
        RECT 393.950 815.720 397.710 816.410 ;
        RECT 398.550 815.720 402.310 816.410 ;
        RECT 403.150 815.720 406.910 816.410 ;
        RECT 407.750 815.720 411.510 816.410 ;
        RECT 412.350 815.720 416.110 816.410 ;
        RECT 416.950 815.720 420.710 816.410 ;
        RECT 421.550 815.720 425.310 816.410 ;
        RECT 426.150 815.720 429.910 816.410 ;
        RECT 430.750 815.720 434.510 816.410 ;
        RECT 435.350 815.720 439.110 816.410 ;
        RECT 439.950 815.720 443.710 816.410 ;
        RECT 444.550 815.720 448.310 816.410 ;
        RECT 449.150 815.720 452.910 816.410 ;
        RECT 453.750 815.720 457.510 816.410 ;
        RECT 458.350 815.720 462.110 816.410 ;
        RECT 462.950 815.720 466.710 816.410 ;
        RECT 467.550 815.720 471.310 816.410 ;
        RECT 472.150 815.720 475.910 816.410 ;
        RECT 476.750 815.720 480.510 816.410 ;
        RECT 481.350 815.720 485.110 816.410 ;
        RECT 485.950 815.720 489.710 816.410 ;
        RECT 490.550 815.720 494.310 816.410 ;
        RECT 495.150 815.720 498.910 816.410 ;
        RECT 499.750 815.720 503.510 816.410 ;
        RECT 504.350 815.720 508.110 816.410 ;
        RECT 508.950 815.720 512.710 816.410 ;
        RECT 513.550 815.720 517.310 816.410 ;
        RECT 518.150 815.720 521.910 816.410 ;
        RECT 522.750 815.720 526.510 816.410 ;
        RECT 527.350 815.720 531.110 816.410 ;
        RECT 531.950 815.720 535.710 816.410 ;
        RECT 536.550 815.720 540.310 816.410 ;
        RECT 541.150 815.720 544.910 816.410 ;
        RECT 545.750 815.720 549.510 816.410 ;
        RECT 550.350 815.720 554.110 816.410 ;
        RECT 554.950 815.720 558.710 816.410 ;
        RECT 559.550 815.720 563.310 816.410 ;
        RECT 564.150 815.720 567.910 816.410 ;
        RECT 568.750 815.720 572.510 816.410 ;
        RECT 573.350 815.720 577.110 816.410 ;
        RECT 577.950 815.720 581.710 816.410 ;
        RECT 582.550 815.720 586.310 816.410 ;
        RECT 587.150 815.720 589.620 816.410 ;
        RECT 1.480 4.280 589.620 815.720 ;
        RECT 2.030 3.670 3.490 4.280 ;
        RECT 4.330 3.670 5.790 4.280 ;
        RECT 6.630 3.670 8.090 4.280 ;
        RECT 8.930 3.670 10.390 4.280 ;
        RECT 11.230 3.670 12.690 4.280 ;
        RECT 13.530 3.670 14.990 4.280 ;
        RECT 15.830 3.670 17.290 4.280 ;
        RECT 18.130 3.670 19.590 4.280 ;
        RECT 20.430 3.670 21.890 4.280 ;
        RECT 22.730 3.670 24.190 4.280 ;
        RECT 25.030 3.670 26.490 4.280 ;
        RECT 27.330 3.670 28.790 4.280 ;
        RECT 29.630 3.670 31.090 4.280 ;
        RECT 31.930 3.670 33.390 4.280 ;
        RECT 34.230 3.670 35.690 4.280 ;
        RECT 36.530 3.670 37.990 4.280 ;
        RECT 38.830 3.670 40.290 4.280 ;
        RECT 41.130 3.670 42.590 4.280 ;
        RECT 43.430 3.670 44.890 4.280 ;
        RECT 45.730 3.670 47.190 4.280 ;
        RECT 48.030 3.670 49.490 4.280 ;
        RECT 50.330 3.670 51.790 4.280 ;
        RECT 52.630 3.670 54.090 4.280 ;
        RECT 54.930 3.670 56.390 4.280 ;
        RECT 57.230 3.670 58.690 4.280 ;
        RECT 59.530 3.670 60.990 4.280 ;
        RECT 61.830 3.670 63.290 4.280 ;
        RECT 64.130 3.670 65.590 4.280 ;
        RECT 66.430 3.670 67.890 4.280 ;
        RECT 68.730 3.670 70.190 4.280 ;
        RECT 71.030 3.670 72.490 4.280 ;
        RECT 73.330 3.670 74.790 4.280 ;
        RECT 75.630 3.670 77.090 4.280 ;
        RECT 77.930 3.670 79.390 4.280 ;
        RECT 80.230 3.670 81.690 4.280 ;
        RECT 82.530 3.670 83.990 4.280 ;
        RECT 84.830 3.670 86.290 4.280 ;
        RECT 87.130 3.670 88.590 4.280 ;
        RECT 89.430 3.670 90.890 4.280 ;
        RECT 91.730 3.670 93.190 4.280 ;
        RECT 94.030 3.670 95.490 4.280 ;
        RECT 96.330 3.670 97.790 4.280 ;
        RECT 98.630 3.670 100.090 4.280 ;
        RECT 100.930 3.670 102.390 4.280 ;
        RECT 103.230 3.670 104.690 4.280 ;
        RECT 105.530 3.670 106.990 4.280 ;
        RECT 107.830 3.670 109.290 4.280 ;
        RECT 110.130 3.670 111.590 4.280 ;
        RECT 112.430 3.670 113.890 4.280 ;
        RECT 114.730 3.670 116.190 4.280 ;
        RECT 117.030 3.670 118.490 4.280 ;
        RECT 119.330 3.670 120.790 4.280 ;
        RECT 121.630 3.670 123.090 4.280 ;
        RECT 123.930 3.670 125.390 4.280 ;
        RECT 126.230 3.670 127.690 4.280 ;
        RECT 128.530 3.670 129.990 4.280 ;
        RECT 130.830 3.670 132.290 4.280 ;
        RECT 133.130 3.670 134.590 4.280 ;
        RECT 135.430 3.670 136.890 4.280 ;
        RECT 137.730 3.670 139.190 4.280 ;
        RECT 140.030 3.670 141.490 4.280 ;
        RECT 142.330 3.670 143.790 4.280 ;
        RECT 144.630 3.670 146.090 4.280 ;
        RECT 146.930 3.670 148.390 4.280 ;
        RECT 149.230 3.670 150.690 4.280 ;
        RECT 151.530 3.670 152.990 4.280 ;
        RECT 153.830 3.670 155.290 4.280 ;
        RECT 156.130 3.670 157.590 4.280 ;
        RECT 158.430 3.670 159.890 4.280 ;
        RECT 160.730 3.670 162.190 4.280 ;
        RECT 163.030 3.670 164.490 4.280 ;
        RECT 165.330 3.670 166.790 4.280 ;
        RECT 167.630 3.670 169.090 4.280 ;
        RECT 169.930 3.670 171.390 4.280 ;
        RECT 172.230 3.670 173.690 4.280 ;
        RECT 174.530 3.670 175.990 4.280 ;
        RECT 176.830 3.670 178.290 4.280 ;
        RECT 179.130 3.670 180.590 4.280 ;
        RECT 181.430 3.670 182.890 4.280 ;
        RECT 183.730 3.670 185.190 4.280 ;
        RECT 186.030 3.670 187.490 4.280 ;
        RECT 188.330 3.670 189.790 4.280 ;
        RECT 190.630 3.670 192.090 4.280 ;
        RECT 192.930 3.670 194.390 4.280 ;
        RECT 195.230 3.670 196.690 4.280 ;
        RECT 197.530 3.670 198.990 4.280 ;
        RECT 199.830 3.670 201.290 4.280 ;
        RECT 202.130 3.670 203.590 4.280 ;
        RECT 204.430 3.670 205.890 4.280 ;
        RECT 206.730 3.670 208.190 4.280 ;
        RECT 209.030 3.670 210.490 4.280 ;
        RECT 211.330 3.670 212.790 4.280 ;
        RECT 213.630 3.670 215.090 4.280 ;
        RECT 215.930 3.670 217.390 4.280 ;
        RECT 218.230 3.670 219.690 4.280 ;
        RECT 220.530 3.670 221.990 4.280 ;
        RECT 222.830 3.670 224.290 4.280 ;
        RECT 225.130 3.670 226.590 4.280 ;
        RECT 227.430 3.670 228.890 4.280 ;
        RECT 229.730 3.670 231.190 4.280 ;
        RECT 232.030 3.670 233.490 4.280 ;
        RECT 234.330 3.670 235.790 4.280 ;
        RECT 236.630 3.670 238.090 4.280 ;
        RECT 238.930 3.670 240.390 4.280 ;
        RECT 241.230 3.670 242.690 4.280 ;
        RECT 243.530 3.670 244.990 4.280 ;
        RECT 245.830 3.670 247.290 4.280 ;
        RECT 248.130 3.670 249.590 4.280 ;
        RECT 250.430 3.670 251.890 4.280 ;
        RECT 252.730 3.670 254.190 4.280 ;
        RECT 255.030 3.670 256.490 4.280 ;
        RECT 257.330 3.670 258.790 4.280 ;
        RECT 259.630 3.670 261.090 4.280 ;
        RECT 261.930 3.670 263.390 4.280 ;
        RECT 264.230 3.670 265.690 4.280 ;
        RECT 266.530 3.670 267.990 4.280 ;
        RECT 268.830 3.670 270.290 4.280 ;
        RECT 271.130 3.670 272.590 4.280 ;
        RECT 273.430 3.670 274.890 4.280 ;
        RECT 275.730 3.670 277.190 4.280 ;
        RECT 278.030 3.670 279.490 4.280 ;
        RECT 280.330 3.670 281.790 4.280 ;
        RECT 282.630 3.670 284.090 4.280 ;
        RECT 284.930 3.670 286.390 4.280 ;
        RECT 287.230 3.670 288.690 4.280 ;
        RECT 289.530 3.670 290.990 4.280 ;
        RECT 291.830 3.670 293.290 4.280 ;
        RECT 294.130 3.670 295.590 4.280 ;
        RECT 296.430 3.670 297.890 4.280 ;
        RECT 298.730 3.670 300.190 4.280 ;
        RECT 301.030 3.670 302.490 4.280 ;
        RECT 303.330 3.670 304.790 4.280 ;
        RECT 305.630 3.670 307.090 4.280 ;
        RECT 307.930 3.670 309.390 4.280 ;
        RECT 310.230 3.670 311.690 4.280 ;
        RECT 312.530 3.670 313.990 4.280 ;
        RECT 314.830 3.670 316.290 4.280 ;
        RECT 317.130 3.670 318.590 4.280 ;
        RECT 319.430 3.670 320.890 4.280 ;
        RECT 321.730 3.670 323.190 4.280 ;
        RECT 324.030 3.670 325.490 4.280 ;
        RECT 326.330 3.670 327.790 4.280 ;
        RECT 328.630 3.670 330.090 4.280 ;
        RECT 330.930 3.670 332.390 4.280 ;
        RECT 333.230 3.670 334.690 4.280 ;
        RECT 335.530 3.670 336.990 4.280 ;
        RECT 337.830 3.670 339.290 4.280 ;
        RECT 340.130 3.670 341.590 4.280 ;
        RECT 342.430 3.670 343.890 4.280 ;
        RECT 344.730 3.670 346.190 4.280 ;
        RECT 347.030 3.670 348.490 4.280 ;
        RECT 349.330 3.670 350.790 4.280 ;
        RECT 351.630 3.670 353.090 4.280 ;
        RECT 353.930 3.670 355.390 4.280 ;
        RECT 356.230 3.670 357.690 4.280 ;
        RECT 358.530 3.670 359.990 4.280 ;
        RECT 360.830 3.670 362.290 4.280 ;
        RECT 363.130 3.670 364.590 4.280 ;
        RECT 365.430 3.670 366.890 4.280 ;
        RECT 367.730 3.670 369.190 4.280 ;
        RECT 370.030 3.670 371.490 4.280 ;
        RECT 372.330 3.670 373.790 4.280 ;
        RECT 374.630 3.670 376.090 4.280 ;
        RECT 376.930 3.670 378.390 4.280 ;
        RECT 379.230 3.670 380.690 4.280 ;
        RECT 381.530 3.670 382.990 4.280 ;
        RECT 383.830 3.670 385.290 4.280 ;
        RECT 386.130 3.670 387.590 4.280 ;
        RECT 388.430 3.670 389.890 4.280 ;
        RECT 390.730 3.670 392.190 4.280 ;
        RECT 393.030 3.670 394.490 4.280 ;
        RECT 395.330 3.670 396.790 4.280 ;
        RECT 397.630 3.670 399.090 4.280 ;
        RECT 399.930 3.670 401.390 4.280 ;
        RECT 402.230 3.670 403.690 4.280 ;
        RECT 404.530 3.670 405.990 4.280 ;
        RECT 406.830 3.670 408.290 4.280 ;
        RECT 409.130 3.670 410.590 4.280 ;
        RECT 411.430 3.670 412.890 4.280 ;
        RECT 413.730 3.670 415.190 4.280 ;
        RECT 416.030 3.670 417.490 4.280 ;
        RECT 418.330 3.670 419.790 4.280 ;
        RECT 420.630 3.670 422.090 4.280 ;
        RECT 422.930 3.670 424.390 4.280 ;
        RECT 425.230 3.670 426.690 4.280 ;
        RECT 427.530 3.670 428.990 4.280 ;
        RECT 429.830 3.670 431.290 4.280 ;
        RECT 432.130 3.670 433.590 4.280 ;
        RECT 434.430 3.670 435.890 4.280 ;
        RECT 436.730 3.670 438.190 4.280 ;
        RECT 439.030 3.670 440.490 4.280 ;
        RECT 441.330 3.670 442.790 4.280 ;
        RECT 443.630 3.670 445.090 4.280 ;
        RECT 445.930 3.670 447.390 4.280 ;
        RECT 448.230 3.670 449.690 4.280 ;
        RECT 450.530 3.670 451.990 4.280 ;
        RECT 452.830 3.670 454.290 4.280 ;
        RECT 455.130 3.670 456.590 4.280 ;
        RECT 457.430 3.670 458.890 4.280 ;
        RECT 459.730 3.670 461.190 4.280 ;
        RECT 462.030 3.670 463.490 4.280 ;
        RECT 464.330 3.670 465.790 4.280 ;
        RECT 466.630 3.670 468.090 4.280 ;
        RECT 468.930 3.670 470.390 4.280 ;
        RECT 471.230 3.670 472.690 4.280 ;
        RECT 473.530 3.670 474.990 4.280 ;
        RECT 475.830 3.670 477.290 4.280 ;
        RECT 478.130 3.670 479.590 4.280 ;
        RECT 480.430 3.670 481.890 4.280 ;
        RECT 482.730 3.670 484.190 4.280 ;
        RECT 485.030 3.670 486.490 4.280 ;
        RECT 487.330 3.670 488.790 4.280 ;
        RECT 489.630 3.670 491.090 4.280 ;
        RECT 491.930 3.670 493.390 4.280 ;
        RECT 494.230 3.670 495.690 4.280 ;
        RECT 496.530 3.670 497.990 4.280 ;
        RECT 498.830 3.670 500.290 4.280 ;
        RECT 501.130 3.670 502.590 4.280 ;
        RECT 503.430 3.670 504.890 4.280 ;
        RECT 505.730 3.670 507.190 4.280 ;
        RECT 508.030 3.670 509.490 4.280 ;
        RECT 510.330 3.670 511.790 4.280 ;
        RECT 512.630 3.670 514.090 4.280 ;
        RECT 514.930 3.670 516.390 4.280 ;
        RECT 517.230 3.670 518.690 4.280 ;
        RECT 519.530 3.670 520.990 4.280 ;
        RECT 521.830 3.670 523.290 4.280 ;
        RECT 524.130 3.670 525.590 4.280 ;
        RECT 526.430 3.670 527.890 4.280 ;
        RECT 528.730 3.670 530.190 4.280 ;
        RECT 531.030 3.670 532.490 4.280 ;
        RECT 533.330 3.670 534.790 4.280 ;
        RECT 535.630 3.670 537.090 4.280 ;
        RECT 537.930 3.670 539.390 4.280 ;
        RECT 540.230 3.670 541.690 4.280 ;
        RECT 542.530 3.670 543.990 4.280 ;
        RECT 544.830 3.670 546.290 4.280 ;
        RECT 547.130 3.670 548.590 4.280 ;
        RECT 549.430 3.670 550.890 4.280 ;
        RECT 551.730 3.670 553.190 4.280 ;
        RECT 554.030 3.670 555.490 4.280 ;
        RECT 556.330 3.670 557.790 4.280 ;
        RECT 558.630 3.670 560.090 4.280 ;
        RECT 560.930 3.670 562.390 4.280 ;
        RECT 563.230 3.670 564.690 4.280 ;
        RECT 565.530 3.670 566.990 4.280 ;
        RECT 567.830 3.670 569.290 4.280 ;
        RECT 570.130 3.670 571.590 4.280 ;
        RECT 572.430 3.670 573.890 4.280 ;
        RECT 574.730 3.670 576.190 4.280 ;
        RECT 577.030 3.670 578.490 4.280 ;
        RECT 579.330 3.670 580.790 4.280 ;
        RECT 581.630 3.670 583.090 4.280 ;
        RECT 583.930 3.670 585.390 4.280 ;
        RECT 586.230 3.670 587.690 4.280 ;
        RECT 588.530 3.670 589.620 4.280 ;
      LAYER met3 ;
        RECT 4.000 808.840 585.600 809.700 ;
        RECT 4.000 800.720 586.000 808.840 ;
        RECT 4.400 799.320 586.000 800.720 ;
        RECT 4.000 793.240 586.000 799.320 ;
        RECT 4.000 791.840 585.600 793.240 ;
        RECT 4.000 776.240 586.000 791.840 ;
        RECT 4.000 774.840 585.600 776.240 ;
        RECT 4.000 772.840 586.000 774.840 ;
        RECT 4.400 771.440 586.000 772.840 ;
        RECT 4.000 759.240 586.000 771.440 ;
        RECT 4.000 757.840 585.600 759.240 ;
        RECT 4.000 744.960 586.000 757.840 ;
        RECT 4.400 743.560 586.000 744.960 ;
        RECT 4.000 742.240 586.000 743.560 ;
        RECT 4.000 740.840 585.600 742.240 ;
        RECT 4.000 725.240 586.000 740.840 ;
        RECT 4.000 723.840 585.600 725.240 ;
        RECT 4.000 717.080 586.000 723.840 ;
        RECT 4.400 715.680 586.000 717.080 ;
        RECT 4.000 708.240 586.000 715.680 ;
        RECT 4.000 706.840 585.600 708.240 ;
        RECT 4.000 691.240 586.000 706.840 ;
        RECT 4.000 689.840 585.600 691.240 ;
        RECT 4.000 689.200 586.000 689.840 ;
        RECT 4.400 687.800 586.000 689.200 ;
        RECT 4.000 674.240 586.000 687.800 ;
        RECT 4.000 672.840 585.600 674.240 ;
        RECT 4.000 661.320 586.000 672.840 ;
        RECT 4.400 659.920 586.000 661.320 ;
        RECT 4.000 657.240 586.000 659.920 ;
        RECT 4.000 655.840 585.600 657.240 ;
        RECT 4.000 640.240 586.000 655.840 ;
        RECT 4.000 638.840 585.600 640.240 ;
        RECT 4.000 633.440 586.000 638.840 ;
        RECT 4.400 632.040 586.000 633.440 ;
        RECT 4.000 623.240 586.000 632.040 ;
        RECT 4.000 621.840 585.600 623.240 ;
        RECT 4.000 606.240 586.000 621.840 ;
        RECT 4.000 605.560 585.600 606.240 ;
        RECT 4.400 604.840 585.600 605.560 ;
        RECT 4.400 604.160 586.000 604.840 ;
        RECT 4.000 589.240 586.000 604.160 ;
        RECT 4.000 587.840 585.600 589.240 ;
        RECT 4.000 577.680 586.000 587.840 ;
        RECT 4.400 576.280 586.000 577.680 ;
        RECT 4.000 572.240 586.000 576.280 ;
        RECT 4.000 570.840 585.600 572.240 ;
        RECT 4.000 555.240 586.000 570.840 ;
        RECT 4.000 553.840 585.600 555.240 ;
        RECT 4.000 549.800 586.000 553.840 ;
        RECT 4.400 548.400 586.000 549.800 ;
        RECT 4.000 538.240 586.000 548.400 ;
        RECT 4.000 536.840 585.600 538.240 ;
        RECT 4.000 521.920 586.000 536.840 ;
        RECT 4.400 521.240 586.000 521.920 ;
        RECT 4.400 520.520 585.600 521.240 ;
        RECT 4.000 519.840 585.600 520.520 ;
        RECT 4.000 504.240 586.000 519.840 ;
        RECT 4.000 502.840 585.600 504.240 ;
        RECT 4.000 494.040 586.000 502.840 ;
        RECT 4.400 492.640 586.000 494.040 ;
        RECT 4.000 487.240 586.000 492.640 ;
        RECT 4.000 485.840 585.600 487.240 ;
        RECT 4.000 470.240 586.000 485.840 ;
        RECT 4.000 468.840 585.600 470.240 ;
        RECT 4.000 466.160 586.000 468.840 ;
        RECT 4.400 464.760 586.000 466.160 ;
        RECT 4.000 453.240 586.000 464.760 ;
        RECT 4.000 451.840 585.600 453.240 ;
        RECT 4.000 438.280 586.000 451.840 ;
        RECT 4.400 436.880 586.000 438.280 ;
        RECT 4.000 436.240 586.000 436.880 ;
        RECT 4.000 434.840 585.600 436.240 ;
        RECT 4.000 419.240 586.000 434.840 ;
        RECT 4.000 417.840 585.600 419.240 ;
        RECT 4.000 410.400 586.000 417.840 ;
        RECT 4.400 409.000 586.000 410.400 ;
        RECT 4.000 402.240 586.000 409.000 ;
        RECT 4.000 400.840 585.600 402.240 ;
        RECT 4.000 385.240 586.000 400.840 ;
        RECT 4.000 383.840 585.600 385.240 ;
        RECT 4.000 382.520 586.000 383.840 ;
        RECT 4.400 381.120 586.000 382.520 ;
        RECT 4.000 368.240 586.000 381.120 ;
        RECT 4.000 366.840 585.600 368.240 ;
        RECT 4.000 354.640 586.000 366.840 ;
        RECT 4.400 353.240 586.000 354.640 ;
        RECT 4.000 351.240 586.000 353.240 ;
        RECT 4.000 349.840 585.600 351.240 ;
        RECT 4.000 334.240 586.000 349.840 ;
        RECT 4.000 332.840 585.600 334.240 ;
        RECT 4.000 326.760 586.000 332.840 ;
        RECT 4.400 325.360 586.000 326.760 ;
        RECT 4.000 317.240 586.000 325.360 ;
        RECT 4.000 315.840 585.600 317.240 ;
        RECT 4.000 300.240 586.000 315.840 ;
        RECT 4.000 298.880 585.600 300.240 ;
        RECT 4.400 298.840 585.600 298.880 ;
        RECT 4.400 297.480 586.000 298.840 ;
        RECT 4.000 283.240 586.000 297.480 ;
        RECT 4.000 281.840 585.600 283.240 ;
        RECT 4.000 271.000 586.000 281.840 ;
        RECT 4.400 269.600 586.000 271.000 ;
        RECT 4.000 266.240 586.000 269.600 ;
        RECT 4.000 264.840 585.600 266.240 ;
        RECT 4.000 249.240 586.000 264.840 ;
        RECT 4.000 247.840 585.600 249.240 ;
        RECT 4.000 243.120 586.000 247.840 ;
        RECT 4.400 241.720 586.000 243.120 ;
        RECT 4.000 232.240 586.000 241.720 ;
        RECT 4.000 230.840 585.600 232.240 ;
        RECT 4.000 215.240 586.000 230.840 ;
        RECT 4.400 213.840 585.600 215.240 ;
        RECT 4.000 198.240 586.000 213.840 ;
        RECT 4.000 196.840 585.600 198.240 ;
        RECT 4.000 187.360 586.000 196.840 ;
        RECT 4.400 185.960 586.000 187.360 ;
        RECT 4.000 181.240 586.000 185.960 ;
        RECT 4.000 179.840 585.600 181.240 ;
        RECT 4.000 164.240 586.000 179.840 ;
        RECT 4.000 162.840 585.600 164.240 ;
        RECT 4.000 159.480 586.000 162.840 ;
        RECT 4.400 158.080 586.000 159.480 ;
        RECT 4.000 147.240 586.000 158.080 ;
        RECT 4.000 145.840 585.600 147.240 ;
        RECT 4.000 131.600 586.000 145.840 ;
        RECT 4.400 130.240 586.000 131.600 ;
        RECT 4.400 130.200 585.600 130.240 ;
        RECT 4.000 128.840 585.600 130.200 ;
        RECT 4.000 113.240 586.000 128.840 ;
        RECT 4.000 111.840 585.600 113.240 ;
        RECT 4.000 103.720 586.000 111.840 ;
        RECT 4.400 102.320 586.000 103.720 ;
        RECT 4.000 96.240 586.000 102.320 ;
        RECT 4.000 94.840 585.600 96.240 ;
        RECT 4.000 79.240 586.000 94.840 ;
        RECT 4.000 77.840 585.600 79.240 ;
        RECT 4.000 75.840 586.000 77.840 ;
        RECT 4.400 74.440 586.000 75.840 ;
        RECT 4.000 62.240 586.000 74.440 ;
        RECT 4.000 60.840 585.600 62.240 ;
        RECT 4.000 47.960 586.000 60.840 ;
        RECT 4.400 46.560 586.000 47.960 ;
        RECT 4.000 45.240 586.000 46.560 ;
        RECT 4.000 43.840 585.600 45.240 ;
        RECT 4.000 28.240 586.000 43.840 ;
        RECT 4.000 26.840 585.600 28.240 ;
        RECT 4.000 20.080 586.000 26.840 ;
        RECT 4.400 18.680 586.000 20.080 ;
        RECT 4.000 11.240 586.000 18.680 ;
        RECT 4.000 9.840 585.600 11.240 ;
        RECT 4.000 9.015 586.000 9.840 ;
      LAYER met4 ;
        RECT 9.495 808.480 580.225 809.705 ;
        RECT 9.495 10.240 20.640 808.480 ;
        RECT 23.040 10.240 97.440 808.480 ;
        RECT 99.840 10.240 174.240 808.480 ;
        RECT 176.640 10.240 251.040 808.480 ;
        RECT 253.440 10.240 327.840 808.480 ;
        RECT 330.240 10.240 404.640 808.480 ;
        RECT 407.040 10.240 481.440 808.480 ;
        RECT 483.840 10.240 558.240 808.480 ;
        RECT 560.640 10.240 580.225 808.480 ;
        RECT 9.495 9.015 580.225 10.240 ;
  END
END RF
END LIBRARY

